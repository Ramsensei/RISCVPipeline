`include "./top/Controller.sv"
`include "./top/IFPipe.sv"
`include "./top/IDPipe.sv"
`include "./top/EXPipe.sv"
`include "./top/MEMPipe.sv"
`include "./top/WBPipe.sv"
`include "./top/IF_IDReg.sv"
`include "./top/ID_EXReg.sv"
`include "./top/EX_MEMReg.sv"
`include "./top/MEM_WBReg.sv"
`define TOP
`include "./components/Mux.sv"
`include "./components/Adder.sv"

module top(clk, rst);

    input clk;
    input rst;

    
    
    
    
endmodule